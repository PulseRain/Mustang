
`timescale 1ns/1ps

parameter CLK_PERIOD =  83.34ns;
parameter unsigned [7 : 0] DEBUG_ADDR = 8'hC0;



module tb_soc ();
    
    logic clk = 0;
    bit reset_n;
    
    logic  start_TX = 0;
    logic  start_RX = 0;
      
    logic unsigned [7 : 0]   data_tx;
    
    wire class_8051_unit_pulse;
       
    wire timer_trigger;
    
    logic test_all_done = 0;
    

    
    int test_case = 0;
    


    
    
    
     Mustang_fast uut (
          
    //=======================================================================
    // clock / reset
    //=======================================================================
            .osc_in (clk),          // expecting 12MHz oscillator in
            .push_button (1'b0),    // push button for reset
        
    //=======================================================================
    // external interrupt
    //=======================================================================
         //   .INTx (2'b00),
    
    //=======================================================================
    // IO port
    //=======================================================================
            .P0 (),
            .P1 (),
     //   inout wire unsigned [7 : 0] P2,
     //   inout wire unsigned [7 : 0] P3,
        
    //=======================================================================
    // UART
    //=======================================================================
            .UART_RXD (1'b0),
            .UART_TXD (),
            
            .UART_AUX_RXD (1'b0),
            .UART_AUX_TXD (),
        
    //=======================================================================
    // debug LED
    //=======================================================================
            .debug_led (),
        
    //=======================================================================
    // M23XX1024
    //=======================================================================
            .mem_so (1'b0),
            .mem_si (),
            .mem_hold_n (),
            .mem_cs_n (),
            .mem_sck (),
          
    //=======================================================================
    // Si3000
    //=======================================================================
            .Si3000_SDO (),
            .Si3000_SDI (),
            .Si3000_SCLK (),
            .Si3000_MCLK (),
            .Si3000_FSYNC_N (1'b0),
            .Si3000_RESET_N (),
          
    //=======================================================================
    // SD Card
    //=======================================================================
            .SD_SPI_CS (),
            .SD_SPI_CLK (),
            .SD_SPI_DO (1'b0),
            .SD_SPI_DI (),
            .SD_DAT2 (),
            .SD_DAT1 (),

    //=======================================================================
    // I2C
    //=======================================================================
            .I2C_SDA (),
            .I2C_SCL (),
        
    //=======================================================================
    // PWM
    //=======================================================================
            .PWM_OUT (),
    //=======================================================================
    // GPIO on JTAG connector
    //=======================================================================
            .JTAG_PIN6 (),
            .JTAG_PIN7 (),
            .JTAG_PIN8 ()
  
);
    
   
    
    initial begin
        forever begin 
            #(CLK_PERIOD/2);
            
            if (test_all_done) begin
                break;
            end else begin
                clk = (~clk);
            end
        end
    end
    
    initial begin
        
        $display ("test start");
        
        
        reset_n = 1;
        # (6 * CLK_PERIOD);
        reset_n = 0;
        
        # (30 * CLK_PERIOD);
        
        reset_n = 1;
        
        # (10 * CLK_PERIOD);
    end            
    
endmodule : tb_soc


